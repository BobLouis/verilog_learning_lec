module test(out1,out2,out3);


	output  [6:0]out1;
	output  [6:0]out2;
    output  [6:0]out3;
		 
	assign out1 = 7'b1000000;
    assign out2 = 7'b1111001;
    assign out3 = 7'b0110000;

endmodule